//
// Table: 0
//
logic [1-1:0][2-1:0][64-1:0][9:0] hash_lup;
// Block: 0
assign hash_lup[0][0][0] = 0;
assign hash_lup[0][0][1] = 134;
assign hash_lup[0][0][2] = 773;
assign hash_lup[0][0][3] = 469;
assign hash_lup[0][0][4] = 545;
assign hash_lup[0][0][5] = 224;
assign hash_lup[0][0][6] = 48;
assign hash_lup[0][0][7] = 695;
assign hash_lup[0][0][8] = 695;
assign hash_lup[0][0][9] = 957;
assign hash_lup[0][0][10] = 392;
assign hash_lup[0][0][11] = 531;
assign hash_lup[0][0][12] = 850;
assign hash_lup[0][0][13] = 35;
assign hash_lup[0][0][14] = 54;
assign hash_lup[0][0][15] = 542;
assign hash_lup[0][0][16] = 687;
assign hash_lup[0][0][17] = 7;
assign hash_lup[0][0][18] = 392;
assign hash_lup[0][0][19] = 68;
assign hash_lup[0][0][20] = 427;
assign hash_lup[0][0][21] = 703;
assign hash_lup[0][0][22] = 603;
assign hash_lup[0][0][23] = 952;
assign hash_lup[0][0][24] = 866;
assign hash_lup[0][0][25] = 539;
assign hash_lup[0][0][26] = 94;
assign hash_lup[0][0][27] = 669;
assign hash_lup[0][0][28] = 425;
assign hash_lup[0][0][29] = 718;
assign hash_lup[0][0][30] = 932;
assign hash_lup[0][0][31] = 780;
assign hash_lup[0][0][32] = 268;
assign hash_lup[0][0][33] = 48;
assign hash_lup[0][0][34] = 753;
assign hash_lup[0][0][35] = 336;
assign hash_lup[0][0][36] = 647;
assign hash_lup[0][0][37] = 774;
assign hash_lup[0][0][38] = 1014;
assign hash_lup[0][0][39] = 374;
assign hash_lup[0][0][40] = 252;
assign hash_lup[0][0][41] = 1006;
assign hash_lup[0][0][42] = 740;
assign hash_lup[0][0][43] = 771;
assign hash_lup[0][0][44] = 667;
assign hash_lup[0][0][45] = 74;
assign hash_lup[0][0][46] = 646;
assign hash_lup[0][0][47] = 905;
assign hash_lup[0][0][48] = 279;
assign hash_lup[0][0][49] = 446;
assign hash_lup[0][0][50] = 784;
assign hash_lup[0][0][51] = 489;
assign hash_lup[0][0][52] = 243;
assign hash_lup[0][0][53] = 281;
assign hash_lup[0][0][54] = 367;
assign hash_lup[0][0][55] = 170;
assign hash_lup[0][0][56] = 498;
assign hash_lup[0][0][57] = 919;
assign hash_lup[0][0][58] = 931;
assign hash_lup[0][0][59] = 62;
assign hash_lup[0][0][60] = 926;
assign hash_lup[0][0][61] = 516;
assign hash_lup[0][0][62] = 528;
assign hash_lup[0][0][63] = 326;

// Block: 1
assign hash_lup[0][1][0] = 1010;
assign hash_lup[0][1][1] = 505;
assign hash_lup[0][1][2] = 272;
assign hash_lup[0][1][3] = 92;
assign hash_lup[0][1][4] = 970;
assign hash_lup[0][1][5] = 75;
assign hash_lup[0][1][6] = 512;
assign hash_lup[0][1][7] = 393;
assign hash_lup[0][1][8] = 283;
assign hash_lup[0][1][9] = 935;
assign hash_lup[0][1][10] = 542;
assign hash_lup[0][1][11] = 475;
assign hash_lup[0][1][12] = 963;
assign hash_lup[0][1][13] = 51;
assign hash_lup[0][1][14] = 779;
assign hash_lup[0][1][15] = 788;
assign hash_lup[0][1][16] = 847;
assign hash_lup[0][1][17] = 128;
assign hash_lup[0][1][18] = 16;
assign hash_lup[0][1][19] = 704;
assign hash_lup[0][1][20] = 889;
assign hash_lup[0][1][21] = 644;
assign hash_lup[0][1][22] = 753;
assign hash_lup[0][1][23] = 742;
assign hash_lup[0][1][24] = 1023;
assign hash_lup[0][1][25] = 909;
assign hash_lup[0][1][26] = 238;
assign hash_lup[0][1][27] = 313;
assign hash_lup[0][1][28] = 359;
assign hash_lup[0][1][29] = 525;
assign hash_lup[0][1][30] = 605;
assign hash_lup[0][1][31] = 866;
assign hash_lup[0][1][32] = 421;
assign hash_lup[0][1][33] = 861;
assign hash_lup[0][1][34] = 275;
assign hash_lup[0][1][35] = 425;
assign hash_lup[0][1][36] = 550;
assign hash_lup[0][1][37] = 479;
assign hash_lup[0][1][38] = 294;
assign hash_lup[0][1][39] = 182;
assign hash_lup[0][1][40] = 157;
assign hash_lup[0][1][41] = 585;
assign hash_lup[0][1][42] = 821;
assign hash_lup[0][1][43] = 33;
assign hash_lup[0][1][44] = 547;
assign hash_lup[0][1][45] = 510;
assign hash_lup[0][1][46] = 978;
assign hash_lup[0][1][47] = 766;
assign hash_lup[0][1][48] = 567;
assign hash_lup[0][1][49] = 912;
assign hash_lup[0][1][50] = 639;
assign hash_lup[0][1][51] = 862;
assign hash_lup[0][1][52] = 163;
assign hash_lup[0][1][53] = 217;
assign hash_lup[0][1][54] = 731;
assign hash_lup[0][1][55] = 133;
assign hash_lup[0][1][56] = 93;
assign hash_lup[0][1][57] = 281;
assign hash_lup[0][1][58] = 3;
assign hash_lup[0][1][59] = 424;
assign hash_lup[0][1][60] = 27;
assign hash_lup[0][1][61] = 726;
assign hash_lup[0][1][62] = 960;
assign hash_lup[0][1][63] = 245;

